** sch_path: /home/thaonguyen06/eda/project/nand_tran.sch
**.subckt nand_tran
X1 VinA VinB VDD GND Vout nand
Vdd VDD GND 1.8
.save i(vdd)
Vin2 VinA GND pulse(0 1.8 1ns 1ns 1ns 4ns 10ns)
.save i(vin2)
Vin1 VinB GND pulse(0 1.8 10ns 1ns 1ns 4ns 10ns)
.save i(vin1)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran 0.01n 1u
.save all

**** end user architecture code
**.ends

* expanding   symbol:  nand.sym # of pins=5
** sym_path: /home/thaonguyen06/eda/project/nand.sym
** sch_path: /home/thaonguyen06/eda/project/nand.sch
.subckt nand A B VP VN Y
*.opin Y
*.iopin VP
*.iopin VN
*.ipin A
*.ipin B
XM5 Y B net1 VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 A VN net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y B VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
