** sch_path: /home/thaonguyen06/eda/project/celltests/buffer_tran.sch
**.subckt buffer_tran
X1 Vin Vout VDD GND buffer
Vdd VDD GND 1.8
.save i(vdd)
Vin Vin GND pulse(0 1.8 1ns 1ns 1ns 4ns 10ns)
.save i(vin)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/thaonguyen06/eda/uniccass/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


.tran 0.01n 1u
.save all

**** end user architecture code
**.ends

* expanding   symbol:  buffer.sym # of pins=4
** sym_path: /home/thaonguyen06/eda/project/celltests/buffer.sym
** sch_path: /home/thaonguyen06/eda/project/celltests/buffer.sch
.subckt buffer A Y VP VN
*.ipin A
*.iopin VP
*.iopin VN
*.opin Y
X1 A net1 VP VN Inverter
X2 net1 Y VP VN Inverter
.ends


* expanding   symbol:  Inverter.sym # of pins=4
** sym_path: /home/thaonguyen06/eda/project/celltests/Inverter.sym
** sch_path: /home/thaonguyen06/eda/project/celltests/Inverter.sch
.subckt Inverter A Y VP VN
*.ipin A
*.iopin VP
*.opin Y
*.iopin VN
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
